    .INIT_00(256'h01df001d00201101003ff00b002010c000bf392021625000022dfa2020d20b98),
    .INIT_01(256'h01df021d00303fff00b23c0b00220b88001f002021f25000032e0e3280a20b6a),
    .INIT_02(256'h013a00208fa20b9801390020b1203cff0108202022803dfe032e0e3280a03eff),
    .INIT_03(256'h00b2382090c01010001f000100020202022e072090020a56011f010504025000),
    .INIT_04(256'h0139000d080010140108200900d01100032e17220082020601cf502093a01100),
    .INIT_05(256'h001f000d04020202022e100900d20b4c011f012500025000013a003681220b81),
    .INIT_06(256'h0139000150a011000118010144020206032e1f250000110001cf303681601014),
    .INIT_07(256'h02f8100d01020b52022e180b01425000011f010b21520b810138000130001014),
    .INIT_08(256'h014006142002020600b0130d00801100003a03143000101802f9111420020202),
    .INIT_09(256'h037000190012500002fa120110120b81004a0003007010180140061430001100),
    .INIT_0A(256'h00b237102400110000be31228270101c00bd3014106202020250003a82b20b5c),
    .INIT_0B(256'h001f000900820b81001a002d209011000019002d30a0101c0018001235020206),
    .INIT_0C(256'h0129e02df0703eff0108d02081603fff032e372500020b8801cf200201025000),
    .INIT_0D(256'h00bf392dd0705e00022e302081605f00011f012de0703cff013a002081603dfe),
    .INIT_0E(256'h001f002db0725000032e442081620b9801df002dc0705c00003ff02081605d01),
    .INIT_0F(256'h0108200146c01100032e44250000101001df022da072020200b23c2081620a56),
    .INIT_10(256'h022e3d0b01420b81011f010b21501014013a0001300011000139000150020231),
    .INIT_11(256'h01cf000d0080101400b037143002020200b2381420020b4c001f000d01025000),
    .INIT_12(256'h013a00011010101401390003007011000108201430020231032e4e1420001100),
    .INIT_13(256'h00b2032284c20202001f001410620b52022e463a85025000011f011900120b81),
    .INIT_14(256'h0139002d209011000108202d30a20231032e57123500110001cf501024001018),
    .INIT_15(256'h001f002d20920b5c022e502d30a25000011f010601020b81013a000900801018),
    .INIT_16(256'h01390014b002023101180114a0601100032e5f250000101c01cf302d00820202),
    .INIT_17(256'h02f81014f0025000022e5814e0020b81011f0114d000110001380014c000101c),
    .INIT_18(256'h01400614d080901100b01314e082f01e003a0314f0e2f03202f9112500001000),
    .INIT_19(256'h037000250001d00802fa1214a0809012004a0014b083229301400614c080d008),
    .INIT_1A(256'h02f503390001d002009508190e932278020e7d390001d004025000110b93226f),
    .INIT_1B(256'h02f605390000100002f504110073228a0096083e8721d0010095081901132281),
    .INIT_1C(256'h02f63125000362ed02f5301100a0d040009608250000900f009508190f62f001),
    .INIT_1D(256'h02f638208ef362d702f537208860d0800096082087c362ed00950800c000d020),
    .INIT_1E(256'h02f606250000d00802f53c208ef0900f009608208862f0010095082087c01001),
    .INIT_1F(256'h00110014c060d01000160714100362ed0015ef14c060d00402500001100362ed),
    .INIT_20(256'h02500014c060901002d10b141002f00102d60a14c060100202d50914100362d7),
    .INIT_21(256'h00b9113a889362ed00b8101d10a0d020020e6925000362ed037001141000d040),
    .INIT_22(256'h02fa3601a002f00102f935250000100302f83411130362d700ba12111070d080),
    .INIT_23(256'h00b431390000d00400b33020868362ed00bd37090060d008001200208f209010),
    .INIT_24(256'h03ae9b368910900e01ba0019101362d701a9402085a0d01001883001104362ed),
    .INIT_25(256'h02fa36208ef362d002f935208860d04002f83400100362d301120104a000d080),
    .INIT_26(256'h00b8340110d362ca022e90250000d010032ec73688c362cd01c2d0192010d020),
    .INIT_27(256'h0012000115f0901602f20f228ef322a600ba36011200d00400b935228ef0900e),
    .INIT_28(256'h032f59011311d00e01d401228ef0300f0094080113e2b04e001300228ef2f033),
    .INIT_29(256'h03aeae011300d02001ba00228ef0900d01b90001133222b9018840228ef362b8),
    .INIT_2A(256'h02f93501132362ad02f834228ef1d0490133000113109006011201228ef362b8),
    .INIT_2B(256'h00b93501134208df00b834228ef362b8022ea1011331d05302fa36228ef222b9),
    .INIT_2C(256'h02f80c011362094302f20d228ef0130002f30e011350b20200ba36228ef2089b),
    .INIT_2D(256'h00b70f011382093a00b60e228ef362b300b50d011371c32000b40c228ef11301),
    .INIT_2E(256'h014700011412020d014608228ef2089b01460801139208cb00b30e228ef22008),
    .INIT_2F(256'h00b01301143322c502f70e228ef1d002014700011420b002014308228ef20216),
    .INIT_30(256'h01400601145322c5014006228ef1d003014006011440b002014006228ef2021f),
    .INIT_31(256'h00b439011472090c025000228ef010000370000114620b1202f00f228ef20228),
    .INIT_32(256'h00b43c0114901080032efd228ef2b10e01d40001148220080034f0228ef2093a),
    .INIT_33(256'h01ba000114b222eb01b900228ef010400188400114a2b20e001200228ef222eb),
    .INIT_34(256'h02f9350114d20b3e02f834228ef222eb0112010114c0102003aed8228ef2b40e),
    .INIT_35(256'h022ecd0114f20b3e032efd228ef222eb01d2020114e0101002fa36228ef2b80e),
    .INIT_36(256'h02f20f011511d00100ba36228ef322e100b935011501d00000b834228ef0b001),
    .INIT_37(256'h01b900011531d003018840228ef322e5019402011521d00200b43c228ef322e3),
    .INIT_38(256'h00b935011552b10f00b834228ef222ea03ef59011542b80f01ba00228ef322e8),
    .INIT_39(256'h00330101157222ea000380228ef2d01000b20f011560108000ba36228ef222ea),
    .INIT_3A(256'h02f80d011592f01e02f30c228ef01008014808011582d01001490e228ef01010),
    .INIT_3B(256'h014200208f60b002014908228ef202160149080115a2020d000390228ef223ec),
    .INIT_3C(256'h0013020d0200b00202f20e0900d2021f01420625000322f70143082d1061d002),
    .INIT_3D(256'h0140060d0100b0010140060900d2022801400625000322f700b013368f21d003),
    .INIT_3E(256'h037000030603230302f30f090001d0010043002500032300014006368f61d000),
    .INIT_3F(256'h018840250003230b0012000309f1d00300b4380900032306025000250001d002),
    .INIT_40(256'h011201041002b08f03af0a208fd2230f01ba00031602b20f01b900001002b40f),
    .INIT_41(256'h01c2d02089d2d01002fa36208bf0104002f935208c52230f02f8342d1002b04f),
    .INIT_42(256'h00b935250000100800b8342089b2230f022eff208742d010032f2c208fa01020),
    .INIT_43(256'h019402041000100100b438208fa2d01002f20f0319f0100400ba36001002d010),
    .INIT_44(256'h03ef592089d0b23701ba00208bf1980101b900208df0982f0188402d1002f01e),
    .INIT_45(256'h00b20f208fd1d00100ba36329363231d00b9351d0011d00000b8340b0320b001),
    .INIT_46(256'h000390208df1d00302f80d250003233602f30c2089b1d0020013002087432328),
    .INIT_47(256'h0143082087420b6a01420001002011020149082089d010a0014908208bf32346),
    .INIT_48(256'h00b0130319f2fd0d001303001002fc0c02f20e2500003f070142002089b20b95),
    .INIT_49(256'h01400625000223580140062d10020b9b014006041002ff0f014006208fa2fe0e),
    .INIT_4A(256'h0250002d103010a00370000b13220a5602f30f2092220b0c0043000100020a56),
    .INIT_4B(256'h01b9000b03203f070188402089d20b95001200208bf20b6a00b403208df01102),
    .INIT_4C(256'h02f834208742ff0f011201010402fe0e03af37329362fd0d01ba001d0012fc0c),
    .INIT_4D(256'h00b8342087420b0c022f2e0102020a5602fa36250002235b02f9352089b20b9e),
    .INIT_4E(256'h00b4031d000010a002f20f208fd20a5600ba362500020b0c00b9352089b20a56),
    .INIT_4F(256'h01ba002089d03f0701b900208a120b95018840208d720b6a0194023294101102),
    .INIT_50(256'h00ba36208df2ff0f00b9352293e2fe0e00b834208cb2fd0d03ef59250002fc0c),
    .INIT_51(256'h02f80d2087520b0c02f30c00c3020a560013002089d2235e00b20f208d520ba1),
    .INIT_52(256'h014200208dd20b0c0149082090520a560149082091120b0c0003902089b20a56),
    .INIT_53(256'h0013042087520b6a02f20e0bc3a011020142002089d010a0014308208cb20a56),
    .INIT_54(256'h014006208c52fd0d014006208d32fc0c0140062500003f0700b0132089b20b95),
    .INIT_55(256'h0370000bc062236102f30f208a720ba4004300208a72ff0f0140062089d2fe0e),
    .INIT_56(256'h02f20d0bc0420a8b02f20c20875223630012ff0bc0520bef0250002087520a84),
    .INIT_57(256'h025000208e120bef037000209a820a9502f20f2089b2236302f20e2087520bef),
    .INIT_58(256'h020f7d0d5040b01600b1170950220bef00b0162089d20aa1001300208bd22363),
    .INIT_59(256'h00130109c1c0b01802f2202297e1f00002f117209ba0b01702f0163a9671d000),
    .INIT_5A(256'h02f0180bb130b01a020f7d09f1f1f00000b11909e1e0b01900b01809d1d1f000),
    .INIT_5B(256'h00b01a13d000b01c00130210cb01f00002f22114b060b01b02f11914b061f000),
    .INIT_5C(256'h02f11b2fe363639802f01a2ff3b1f000020f7d13f000b01d00b11b13e001f000),
    .INIT_5D(256'h00b11d208752023c00b01c0bc3b2f03a0013032fc341100102f2222fd350b03a),
    .INIT_5E(256'h02f223208753238102f11d0bc351d00202f01c208750b002020f7d0bc3620245),
    .INIT_5F(256'h01f1ff208bf3238101d0ff2089b1d003001200208750b0020250000bc342024e),
    .INIT_60(256'h0140063a9862b08f0140060d5042b20f0140062089d2b40f031000208bd20257),
    .INIT_61(256'h0141000bd35010200140060bc342d0100141002299c01040014006209ba2b04f),
    .INIT_62(256'h01003001b000100401400e01a042d01001400e0bf3b0100801400e0be362d010),
    .INIT_63(256'h022ffc2081201080022ffc09f072b10f025000208122b80f00b224208322d010),
    .INIT_64(256'h022ffc2081220b12022ffc09d072d010022ffc2081201010022ffc09e072d010),
    .INIT_65(256'h022ffc2087522008022ffc00cd0326cf022ffc208751d001022ffc09c070b032),
    .INIT_66(256'h022ffc208752f034022ffc00cf00b016022ffc20875323e7022ffc00ce01d800),
    .INIT_67(256'h022ffc2089d2f036022ffc208d10b018022ffc208bf2f035022ffc2089b0b017),
    .INIT_68(256'h022ffc14c002f03c022ffc0d5040b01a022ffc01c002f03b022ffc208a70b019),
    .INIT_69(256'h022ffc250002f03e022ffc2089b0b01c022ffc208752f03d022ffc11c010b01b),
    .INIT_6A(256'h022ffc2b80c1d000022ffc2089d0b001022ffc208df2f03f022ffc208e10b01d),
    .INIT_6B(256'h022ffc2b02c1d002022ffc20875323b7022ffc09c0c1d001022ffc2b03c323b3),
    .INIT_6C(256'h022ffc09c0c20b9b022ffc2b01c323bf022ffc208751d003022ffc09c0c323bb),
    .INIT_6D(256'h022ffc2087520b9e022ffc09c0c223c2022ffc2b00c20bef022ffc2087520a84),
    .INIT_6E(256'h022ffc208e920ba1022ffc208e9223c2022ffc2500020bef022ffc2089b20a8b),
    .INIT_6F(256'h022ffc208e920ba4022ffc208e9223c2022ffc208e920bef022ffc208e920a95),
    .INIT_70(256'h022ffc0b0320b134022ffc250000b016022ffc208e920bef022ffc208e920aa1),
    .INIT_71(256'h022ffc208d71e010022ffc208bf0b135022ffc369ca0b017022ffc1d0001c010),
    .INIT_72(256'h022ffc208bf0b019022ffc250001e010022ffc2089b0b136022ffc208dd0b018),
    .INIT_73(256'h022ffc250000b13c022ffc2089b0b01a022ffc208bb1e010022ffc208d10b13b),
    .INIT_74(256'h022ffc208c31e010022ffc369d70b13d022ffc1d0000b01b022ffc0b0321e010),
    .INIT_75(256'h022ffc250000b01d022ffc2089b1e010022ffc208c10b13e022ffc208d50b01c),
    .INIT_76(256'h022ffc2089b19801022ffc208bf363fb022ffc208bf1e010022ffc208c30b13f),
    .INIT_77(256'h022ffc2089d1d000022ffc208bb0b001022ffc208d9323e7022ffc209a81d800),
    .INIT_78(256'h022ffc141061d002022ffc14106323b7022ffc141061d001022ffc0b113323b3),
    .INIT_79(256'h022ffc208740b001022ffc04010323bf022ffc0b00f1d003022ffc14106323bb),
    .INIT_7A(256'h022ffc208742f01f022ffc0b00d01004022ffc2087420d8f022ffc0b00e2f013),
    .INIT_7B(256'h022ffc208d11d002022ffc2089b0b032022ffc208742f013022ffc0b00c0b001),
    .INIT_7C(256'h022ffc208740b032022ffc010002094b022ffc2089d2089b022ffc208bb323f2),
    .INIT_7D(256'h022ffc0b0123271b022ffc141061d002022ffc141063271b022ffc0b1131d001),
    .INIT_7E(256'h022ffc208740b03a022ffc0b01122008022ffc208742090c022ffc0401001004),
    .INIT_7F(256'h022ffc250001d00002d0032089b0b0160010ff208742f03a02bff00b01011001),
    .INITP_00(256'h74f1b43f8da8eb932e6c94952eb86787878c481933a129d72a35b04303a42f5b),
    .INITP_01(256'h13c4b09f1269858a0cc989bbba39fc232d8d25a0999030e169503199bf33836e),
    .INITP_02(256'hdb5d9a998f095b3e9ad8b2b6812175048013ff91b9b82d4614899d9c4023050d),
    .INITP_03(256'h90b28d44f3598d03e1521a23c95e148e42f98188de976df564d29e0bb1379764),
    .INITP_04(256'hb5c63390a77bda35d1666aa7ea1dac23371fba1ef0676115a903c352cfd6eb4d),
    .INITP_05(256'h2f7e9b12908d333881b49db9787ee5813b8beefec37dacad6abf8eb0cba99d18),
    .INITP_06(256'hb2a413adc691131c4e692be9ed712f733baca43b38e5058ea8eb6f733ebe2b2a),
    .INITP_07(256'hbc33aae5e2dd01232e0139af2e4f0113a4901bbff5622119840a3f86990e64ac),
    .INITP_08(256'h8f9c048d9ee0e31e880bbd9d622e073fa836e5139a9f656f94715e6d91619ca3),
    .INITP_09(256'h35238238047b1b0e07c7677f72167399a8262c127951ff1ca3a9040e03807095),
    .INITP_0A(256'h44c5cb6dee52b4e9e079152d8a1dbdba2f758323329b14a97b42980ca734267c),
    .INITP_0B(256'ha3b63eea64ccc86426a4126bea5bec859019de6ec052178690e4fe51730cab86),
    .INITP_0C(256'hcc614e41c869c67d597b5cf7f0cbe24ce7ebdd992a0598b82fb510802e37a56c),
    .INITP_0D(256'he2e2e86fe7e2db59de7cf1d8f879d9e6e1447fe75d4c72e5c4404cff62d7c745),
    .INITP_0E(256'h5ed4fa6b5f5fd2634bd17bfb736de5c44f43cee0465945e0f1406de7d54ae8ea),
    .INITP_0F(256'h5152034cd5d44a5540504669d2505953fbced845595c4fd1d7d8d0cf504e56f7),
