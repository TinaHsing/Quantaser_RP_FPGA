    .INIT_00(256'h0000000bc161f00000000034a3e0b0180000001dcff1f0000000000bc170b017),
    .INIT_01(256'h0000001dcff1f0000000000bc190b01a00000034a441f0000000001dcff0b019),
    .INIT_02(256'h00000034a441f0000000001dcff0b01c0000000bc181f00000000034a3e0b01b),
    .INIT_03(256'h0000000bc1a2023c00000034a3e360170000001dcff1f0000000000bc1b0b01d),
    .INIT_04(256'h0000001dcff323810000000bc1d1d00200000034a440b0020000001dcff20245),
    .INIT_05(256'h00000034a44323810000001dcff1d0030000000bc1c0b00200000034a3e2024e),
    .INIT_06(256'h00000032a222b08f0000001dd002b20f0000000bd202b40f0000002500020257),
    .INIT_07(256'h00000020a4a010200000000bc162d01000000020a3e010400000000bc172b04f),
    .INIT_08(256'h0000001dd00010040000000bd212d01000000020a50010080000000bc202d010),
    .INIT_09(256'h0000000bc180108000000020a3e2b10f0000000bc192b80f00000032a2b2d010),
    .INIT_0A(256'h0000000bd2220b1200000020a502d0100000000bc210101000000020a4a2d010),
    .INIT_0B(256'h00000020a3e220080000000bc1b326cf00000032a341d0010000001dd000b032),
    .INIT_0C(256'h00000020a500be110000000bc220bd1000000020a4a2f01e0000000bc1a01001),
    .INIT_0D(256'h0000000bc1d13f0000000032a3d13e000000001dd0011d010000000bd230bf12),
    .INIT_0E(256'h0000000bc232ff1200000020a4a03f030000000bc1c2fe1100000020a3e2fd10),
    .INIT_0F(256'h000000208c12f00f000000208e703007000000250000b00f00000020a5020e84),
    .INIT_10(256'h0000002500003efc0000002089d0be0e00000020875030fc0000002089d0b03b),
    .INIT_11(256'h000000208751d0000000002089d0b001000000208e136477000000208bd1c0e0),
    .INIT_12(256'h000000208e11d002000000208bd32453000000250001d0010000002089b3244f),
    .INIT_13(256'h0000002500020b9b0000002089d3245b000000208751d0030000002089d32457),
    .INIT_14(256'h0000002087520b9e0000002089d2245e000000208e520bef000000208d120a84),
    .INIT_15(256'h0000002b21a20ba10000002bec92245e0000002500020bef0000002089b20a8b),
    .INIT_16(256'h0000002005c20ba400000020bdb2245e0000002b08e20bef0000002b1bb20a95),
    .INIT_17(256'h000000250001d00000000020a6f0b01600000001c0020bef0000002500020aa1),
    .INIT_18(256'h00000001c071f000000000250000b01800000020a6f1f00000000001c100b017),
    .INIT_19(256'h00000020a6f1f00000000001c0d0b01a000000250001f00000000020a6f0b019),
    .INIT_1A(256'h000000250001f00000000020a6f0b01c00000001c011f000000000250000b01b),
    .INIT_1B(256'h00000001d0022477000000250003647000000020a6f1f00000000001c040b01d),
    .INIT_1C(256'h000000010802094b00000020b732089b00000001f002093a00000001e002091b),
    .INIT_1D(256'h000000250002023c00000020a7e2200800000020b6a2090c0000000110001004),
    .INIT_1E(256'h0000002b08e324810000002b63b1d0020000002b00a0b0020000002b38920245),
    .INIT_1F(256'h0000002b00a324810000002b2091d003000000250000b00200000020bdb2024e),
    .INIT_20(256'h000000250002b08f00000020bdb2b20f0000002b08e2b40f0000002b37b20257),
    .INIT_21(256'h0000002b5bb010200000002b62a2d0100000002b6490104000000020a6c2b04f),
    .INIT_22(256'h00000020a5601004000000250002d01000000020bdb010080000002b08e2d010),
    .INIT_23(256'h0000002b6490108000000020a6c2b10f00000020a562b80f00000020b0c2d010),
    .INIT_24(256'h00000020bdb20b120000002b08e2d0100000002b5bb010100000002b62a2d010),
    .INIT_25(256'h00000020a562d01000000020b0c0108000000020a562b10f000000250002b80f),
    .INIT_26(256'h0000002b6492090c00000020a6c0100200000020a562d01000000020b0c01010),
    .INIT_27(256'h00000020bdb2f0320000002b08e010000000002b5bb220080000002b62a2093a),
    .INIT_28(256'h00000020a560901700000020b0c324cd00000020a560d004000000250000900e),
    .INIT_29(256'h00000020a560901900000020b0c2f00800000020a560901800000020b0c2f007),
    .INIT_2A(256'h0000002b5bb0901b0000002b62a2f00a0000002b6490901a00000020a6c2f009),
    .INIT_2B(256'h00000020a692b04e000000250002f03300000020bdb090160000002b08e2f00b),
    .INIT_2C(256'h0000002b08e090020000002bdfb364b70000002b10a1d00a0000002b6490300f),
    .INIT_2D(256'h0000002bebb1d00e0000002b10a226260000002b6c93262500000020bdb0d002),
    .INIT_2E(256'h00000020a56364c4000000250001d00b00000020bdb226250000002b08e364ba),
    .INIT_2F(256'h00000020a56208dd00000020b002dc0100000020b8f03c0f00000001ccc0bc07),
    .INIT_30(256'h0000002bdfb220030000002b10a2089b0000002b6492087500000020a692089d),
    .INIT_31(256'h0000002b10a226370000002b6c9208c100000020bdb364c80000002b08e1d00f),
    .INIT_32(256'h000000250003264c00000020bdb0d0080000002b08e3264c0000002bebb1d00c),
    .INIT_33(256'h00000020b003662500000020b8f0d02000000001cd80900d00000020a5622623),
    .INIT_34(256'h00000020b000900200000020b8f364d700000001ccc1d04f00000020a5609006),
    .INIT_35(256'h0000002b10a1d0530000002b6492262600000020a693262500000020a560d002),
    .INIT_36(256'h0000002b6c90b20200000020bdb2089b0000002b08e208df0000002bdfb364e3),
    .INIT_37(256'h00000020bdb113010000002b08e209520000002bebb209430000002b10a01300),
    .INIT_38(256'h00000020b8f1d05200000001ce42262400000020a56364dd000000250001c320),
    .INIT_39(256'h00000020b8f0900600000001cd8208f200000020a56208dd00000020b00364fa),
    .INIT_3A(256'h00000020b8f208f200000001ccc2089d00000020a563662300000020b001d020),
    .INIT_3B(256'h0000002b649208a700000020a693662300000020a561d03000000020b0009006),
    .INIT_3C(256'h00000020bdb3a6230000002b08e208680000002bdfb090060000002b10a208f2),
    .INIT_3D(256'h0000002b08e208ef0000002bebb208860000002b10a001000000002b6c92d001),
    .INIT_3E(256'h0000002b22a364fe0000002b1c91d044000000250002200300000020bdb2089b),
    .INIT_3F(256'h000000250003652500000020bdb1d04e0000002b08e226370000002b47b208c1),
    .INIT_40(256'h0000002b08e1d0200000002b57b090060000002b22a208f20000002b489208d5),
    .INIT_41(256'h0000002b66a2088b0000002b5c90120a000000250002089d00000020bdb36623),
    .INIT_42(256'h000000250002fc0a00000020bdb2fb090000002b08e2fa080000002b6bb3a623),
    .INIT_43(256'h0000002b08e2088b0000002b7bb012010000002b66a2fe330000002b6c92fd0b),
    .INIT_44(256'h00000020b0c14a0600000020a5614a060000002500014a0600000020bdb3a623),
    .INIT_45(256'h00000020b6a0bd0a000000011010bc09000000010800bb0800000020a5614a06),
    .INIT_46(256'h00000001c0e2086100000020a5620861000000250000bf3300000020a780be0b),
    .INIT_47(256'h00000020a5d2fb0800000020a562fa0700000020b002086100000020b8f20861),
    .INIT_48(256'h00000020b8f2ff3300000001c1e2fe0b00000020a562fd0a000000250002fc09),
    .INIT_49(256'h00000001c0e208e100000020a5d3659200000020a561d05400000020b002265d),
    .INIT_4A(256'h00000020a5d3662300000020a561d02000000020b000900600000020b8f208f2),
    .INIT_4B(256'h00000020b8f3a62300000001c2e2088b00000020a560120a000000250002089d),
    .INIT_4C(256'h00000001c1e2fd0b00000020a5d2fc0a00000020a562fb0900000020b002fa08),
    .INIT_4D(256'h00000020a5d3a62300000020a562088b00000020b000120100000020b8f2fe33),
    .INIT_4E(256'h00000020a5614a0600000020b0014a0600000020b8f14a0600000001c0e3a623),
    .INIT_4F(256'h0000001d0020bb080000000b0020ba07000000250002fa0700000020a5d14a06),
    .INIT_50(256'h0000001d0040bf3300000032b470be0b0000001d0030bd0a00000032b450bc09),
    .INIT_51(256'h00000020b212086100000022b4a2086100000020b1a2086100000032b4920861),
    .INIT_52(256'h000000250002fd0a0000000b0022fc0900000020b2d2fb0800000022b4a2fa07),
    .INIT_53(256'h00000020b002fb3f00000020b8f2fa3e00000001c0e2ff3300000020a562fe0b),
    .INIT_54(256'h00000001c1a3255500000020a560df08000000250003257400000020a561df0c),
    .INIT_55(256'h00000001c0e2085a00000020a562fa1300000020b000ba3300000020b8f22623),
    .INIT_56(256'h000000250002fc0c00000020a562085a00000020b002085a00000020b8f2085a),
    .INIT_57(256'h00000020b0020d8f00000020b8f2ff0f00000001c262fe0e00000020a562fd0d),
    .INIT_58(256'h00000020b000bf1200000020b8f0be1100000001c1a0bd1000000020a562089b),
    .INIT_59(256'h00000020b002087500000020b8f00cf000000001c0e208a700000020a56208bf),
    .INIT_5A(256'h0000002b419208750000002b00a00cd0000000250002087500000020a5600ce0),
    .INIT_5B(256'h0000002b259208860000002b00a2087c0000002d1082087c0000002d0080bc3f),
    .INIT_5C(256'h0000002b00a2262300000025000208750000002d1080bc3e0000002d008208ef),
    .INIT_5D(256'h0000002de082085a0000002dd082fe130000002dc082085a0000002b2892085a),
    .INIT_5E(256'h0000002b2892fd110000002b00a2fc100000002500003e030000002df082085a),
    .INIT_5F(256'h00000009f080bf0c00000009e082089b00000009d0820e8400000009c082fe12),
    .INIT_60(256'h0000002dc08208750000002d0090bc0f0000002d10a0bd0e000000250000be0d),
    .INIT_61(256'h00000025000208750000002df0800ce00000002de08208750000002dd0800cd0),
    .INIT_62(256'h00000009d082087c00000009c080bc3f0000002d009208750000002d10a00cf0),
    .INIT_63(256'h000000010500bc3e00000025000208ef00000009f082088600000009e082087c),
    .INIT_64(256'h0000002dc08365b00000002d0091d0580000002d10a226230000000110220875),
    .INIT_65(256'h00000025000208e900000020b7a3e5b000000020a780d0040000002500009002),
    .INIT_66(256'h00000020a5636623000000250001d02000000020a7e0900600000020b73208f2),
    .INIT_67(256'h00000020ba73a62300000020b4c2088b000000250000120800000020ba72089d),
    .INIT_68(256'h000000250002fc3600000020ba72fb3500000020b522fa34000000250002089b),
    .INIT_69(256'h000000010200be36000000250000bd3500000020ba70bc3400000020b5c2fd3b),
    .INIT_6A(256'h0000000be0e208320000000bf0f01b0000000020b6a01a01000000011000bf3b),
    .INIT_6B(256'h000000250002262300000020b98208750000000bc0c09c070000000bd0d20812),
    .INIT_6C(256'h00000020b6a208f200000001101208db000000010803662500000020b9b1d051),
    .INIT_6D(256'h00000020b982089d00000020b8836623000000011001d0200000000100009006),
    .INIT_6E(256'h00000020b4c2fa0800000020b9e3a623000000250002088b00000020aaf0120a),
    .INIT_6F(256'h000000010042fe3300000020b6a2fd0b000000011012fc0a000000010802fb09),
    .INIT_70(256'h00000020abb14a0600000020b983a62300000020b882088b0000000110001201),
    .INIT_71(256'h000000010800bb0800000020b5214a0600000020ba114a060000002500014a06),
    .INIT_72(256'h000000011000bf33000000010080be0b00000020b6a0bd0a000000011010bc09),
    .INIT_73(256'h000000250002086100000020acc2086100000020b982086100000020b8820861),
    .INIT_74(256'h000000011012fd0a000000010802fc0900000020b5c2fb0800000020ba42fa07),
    .INIT_75(256'h00000020b88325e5000000011001df0c0000000100c2ff3300000020b6a2fe0b),
    .INIT_76(256'h0000000900e2ff13000000250002262300000020ae1325db00000020b980df08),
    .INIT_77(256'h0000000900e2085a000000250002085a00000036bdb2085a0000000d0082085a),
    .INIT_78(256'h0000000900f2ff0f000000250002fe0e00000032bdf2fd0d0000000d0022fc0c),
    .INIT_79(256'h000000090102fe13000000250002085a00000032be32085a0000000d002225fa),
    .INIT_7A(256'h000000090112fc100000002500003e0300000032be72085a0000000d0022085a),
    .INIT_7B(256'h000000370010b105000000250000b00400000032beb2fe120000000d0022fd11),
    .INIT_7C(256'h0000002f1181ae200000002f1171ad100000002f11618c00000000011000b206),
    .INIT_7D(256'h0000002f11c034070000002f11b0b40f0000002f11a20e840000002f1193e623),
    .INIT_7E(256'h0000002b00a0b0130000002b6c920b3e000000010a2225fa0000002f11d2f40f),
    .INIT_7F(256'h00000020c0a3260700000020c051d00100000011001326040000002b00b1d000),
    .INITP_00(256'h1132acaa21a511390f8d282110a38019a5b898bb871233ab98a0871729ad98b8),
    .INITP_01(256'h038ab11c3e93b438a9303b1e1fac13afb6b7b63d889c38043bbc2aa33b0d0434),
    .INITP_02(256'ha70e2b2f17813e1db5a72daf28209f8fa3332fb28c2b24bb29ba0d28362da83b),
    .INITP_03(256'h1d29b39aa3951e3cb917bf90042ea983042306a7b48ca8be06a0b4892fb806a7),
    .INITP_04(256'h1d23b31b24861b171b129fb705bc2b9cb018030102af99bc289c371eaa86ba29),
    .INITP_05(256'h1c94372c9ea6863590a0909ab331aba89b3001273f8422829c9c1f1b98948321),
    .INITP_06(256'h08bd97bd130e3e35ad220b808f28af9285b6219f3b182815aa0e0533352ea596),
    .INITP_07(256'ha9063712bd26200e3d18210b8631332b2e9c100928271d02aba31c022dad93bc),
    .INITP_08(256'h089e892bba122e96309004081208bc863a8bb289a98dbe3dbb95a3073eb7b304),
    .INITP_09(256'h95352a1408933134809d92ada5019782a52a08a301990928360e1708a0a610af),
    .INITP_0A(256'h0222bf90aa108b29b89183a6ab1f3c8f0c203190a4b30b0a8c8611ac9f378b27),
    .INITP_0B(256'h9cb5bd98060f3597b43d108e86a9bb999c80b91b3e1fa90586b53e1808a13214),
    .INITP_0C(256'h272639ac1d2d102b2db586a01d8f2414152e1d38bf1d0437a982b9251d022e24),
    .INITP_0D(256'h39b09584a221290d2db90b2332970da92b27be9418a1bb0f3c23a2b52baea4a0),
    .INITP_0E(256'h91a4203f922bb725aa1da9b3980831a4a62828b608bf3090043734bc8fa6399b),
    .INITP_0F(256'hbaaf8310140e8199921d16048a8a071d27b005b1093509391ba4153f80219537),
