    .INIT_00(256'h0370003260d20020036bfd1d0032ff0001d0ff3260a01f00020c641d00228000),
    .INIT_01(256'h009e0820b9e2090c009d082260f01001009c0820a842004c02500020b9b20033),
    .INIT_02(256'h032c2020a951d00201d0d020ba1320600250002260f1d001009f0820a8b208fd),
    .INIT_03(256'h020c532089b1d0100001f020aa13249e032c3520ba41d00001d0d12260f32260),
    .INIT_04(256'h020c5309f081d0080001d00125d3271b020c532b6c91d0040001e02b00a32669),
    .INIT_05(256'h02f128208750106000110009c0832430020c5309d081d0820001c009e08327c5),
    .INIT_06(256'h02f12920875208c902f12e00ce02090c02f12c208750109f02f12a00cd020900),
    .INIT_07(256'h0250001920122ffc02f12f2089b2089b02f12d20875208e102f12b00cf0208d1),
    .INIT_08(256'h020c532089b0b0000001e0226243202f020c5320b120d0800001f03661309002),
    .INIT_09(256'h020c532089b011ff0001c0208d7010ff020c53220083602f0001d02093a0d001),
    .INIT_0A(256'h02f42e1d0021b20002f52c0b0021b10002f62a202451900102f7282023c0121f),
    .INIT_0B(256'h0017001d003090010016000b0022f0000015002024e01001001400326323e029),
    .INIT_0C(256'h02f42f010022b00002f52d20b122500002f62b202573202f02f729326320d040),
    .INIT_0D(256'h0001e02089b010ff020c53220082bfff0001f02093a2bf7e022c1f2090c2b00c),
    .INIT_0E(256'h0001c01d0020300f020c530b002090010001d0202452d011020c532023c2d010),
    .INIT_0F(256'h02f1291d0033604200310f0b0020d0200001702024e0900d020c53326422d001),
    .INIT_10(256'h02f12b010000900600310f20b1209006000160202572203d0037f03264209006),
    .INIT_11(256'h02f12d209280900700310f2f03236049000150010010d0800036f02f01e0900d),
    .INIT_12(256'h02f12f226cf2500000310f2089d09007000140208a1090070035f0208c122044),
    .INIT_13(256'h02f12a2087c2089f02f1280bc33208d30011002089d208c30034f0208d5208df),
    .INIT_14(256'h0141000bc0b208dd022c1f208ef208e102f12e20886208d102f12c2087c208e3),
    .INIT_15(256'h0141000bc09208a501450020875208e50141000bc0a2089f01440020875208bb),
    .INIT_16(256'h0141000bc0725000014700208752089b0141000bc08208a3014600208752089f),
    .INIT_17(256'h0141000d00825000014500090023e05d0141002089b190010144002087501019),
    .INIT_18(256'h0250002090c0900d01470001010201b501410020b3e201cf01460032665201c7),
    .INIT_19(256'h020d052093a20a5d00b9292090c20a5600b8280100032063000170220080d001),
    .INIT_1A(256'h00ba250bc0920b95001b000bb0820b6a020d2f0ba0701101020d112200801080),
    .INIT_1B(256'h014a00000f00100000ba260bf3301100014b000be0b36066014a0e0bd0a1dc93),
    .INIT_1C(256'h014a000d0080311e014b0032676001e0014a001d00c20e69014b000300f20b81),
    .INIT_1D(256'h02f2170301f320850062b0000a01d11400b217226ca32079014b00326761d112),
    .INIT_1E(256'h014b002085a1410a014a002085a001e0014b002085a000d0014a002f01422017),
    .INIT_1F(256'h014b003e6ca3208f014a001d05d1d058014b000307f030f8014a00000b014008),
    .INIT_20(256'h014a001d00c3209200ba270300f1d088014b000b0333208f014a002f0151d048),
    .INIT_21(256'h014a00000e01410a014b0032690001e0014a000d008000d0014b003268722017),
    .INIT_22(256'h02fb160b11332092006b202f0131d04800b21603003030f8014b001400e14008),
    .INIT_23(256'h020d053669f0100200b92b2085a2201700b82a366ca320950001601c0101d088),
    .INIT_24(256'h00ba250b1132f002001b002f01301003020d2f0300322097020d110b0332f002),
    .INIT_25(256'h014a002fc0c201b100ba262085a2f002014b00366ca01004014a0e1c01022097),
    .INIT_26(256'h014a0003f072f201014b002ff0f01203014a002fe0e2f239014b002fd0d01220),
    .INIT_27(256'h02f21903e032f0240062b0226ae0100100b219326ca2f03a014b001df0101000),
    .INIT_28(256'h014b000b00420202014a002fe12201e3014b002fd11201da014a002fc10201c1),
    .INIT_29(256'h014b001ad1020b81014a0018c0001010014b000b20601100014a000b10520b95),
    .INIT_2A(256'h014a000b40f201ec00ba2720e8401100014b003e6ca01010014a001ae2020202),
    .INIT_2B(256'h014a001d00020a63014b000b01320b81014a002f40f01010014b000340701100),
    .INIT_2C(256'h02fb181d00220bdf006b20326bc2b02e00b2181d00120a66014b00326b720a60),
    .INIT_2D(256'h020d0520b9b20a5600b92d326c620b3e00b82c1d00320bdf000150326c12b02e),
    .INIT_2E(256'h00ba25226ca01101001b0020bb001080020d2f2083f20a56020d1120a8420b0c),
    .INIT_2F(256'h014a0020bba0100400ba262083f01100014b0020a8b20b95014a0e20b9e20b6a),
    .INIT_30(256'h014a002083f20b4c014b0020a95201da014a0020ba120b4c014b00226ca20b81),
    .INIT_31(256'h02f21b20aa120a560062b020ba420b0c00b21b226ca20a56014b0020bc5201e3),
    .INIT_32(256'h014b000100001014014a0020b1201100014b0020bd020b95014a002083f20202),
    .INIT_33(256'h014b000901120b6a014a002200801101014b002093a010c0014a002090c20b81),
    .INIT_34(256'h014a000d080201ec00ba270900e01100014b003626601014014a000d00820b4c),
    .INIT_35(256'h014a000d02020b4c014b00362d020b81014a000d04001014014b00362d301100),
    .INIT_36(256'h02fb1a0900e20b4c006b20362ca20a6000b21a0d01020b4c014b00362cd20a63),
    .INIT_37(256'h020d052f03320be300b92f090162d00f00b82e326e5010020001400d00420a66),
    .INIT_38(256'h00ba25326f90b002001b001d00e20be3020d2f0300f2d00f020d112b04e01002),
    .INIT_39(256'h014a00366cf20a5600ba260d02020b3e014b000900d3214f014a0e226cf1d002),
    .INIT_3A(256'h014a001d05320a56014b00326f920b0c014a001d04920a56014b000900620b0c),
    .INIT_3B(256'h02f21d0b20220b950062b02089b20b6a00b21d208df01101014b00366cf01080),
    .INIT_3C(256'h014b001c32020b52014a001130120b81014b002094301008014a000130001100),
    .INIT_3D(256'h014b002089d20a56014a00208a1201e3014b00208c120b52014a00366f1201da),
    .INIT_3E(256'h014a002020d20a5600ba272089b20b0c014b00208cb20a56014a00226cf20b0c),
    .INIT_3F(256'h014a003270501018014b001d00201100014a000b00220b95014b002021620202),
    .INIT_40(256'h02fb1c3270520b6a006b201d0030110100b21c0b002010c0014b002021f20b81),
    .INIT_41(256'h00d1ff2020d201ec001b002271401100001a0020b12010180250002022820b52),
    .INIT_42(256'h00d9ff3271120b52014a001d00220b8100d8ff0b00201018014a002021601100),
    .INIT_43(256'h02fb253271120b52014b001d00320a6000daff0b00220b52014a002021f20a63),
    .INIT_44(256'h00d1ff2090020be7001a00010602d01000020020b12010020250002022820a66),
    .INIT_45(256'h014a04010000b002014a042d00320be7014a042f0322d010014a000100001002),
    .INIT_46(256'h014a040b01e20a56014a042200820b3e014a042093a3214f014a042090c1d003),
    .INIT_47(256'h0062b00b41620a56020d220120020b0c0022a03678020a56014a041d00120b0c),
    .INIT_48(256'h000b902f91701101000a802f8160108002500020d5320a5602f2260b51720b0c),
    .INIT_49(256'h014b0020d530100c014a060b51901100014b000b41820b95014a060421020b6a),
    .INIT_4A(256'h014b000b41a20b5c014a0604210201da014b002f91920b5c014a062f81820b81),
    .INIT_4B(256'h0002102f91b20a560250002f81a20b0c014b0020d5320a56014a060b51b201e3),
    .INIT_4C(256'h0032aa20d5320a56001b000b51d20b0c001a000b41c20a560003800421020b0c),
    .INIT_4D(256'h00d3ff0d2020101c014a00042100110000d2ff2f91d20b950033012f81c20202),
    .INIT_4E(256'h000210209d820b6a014b082f21e0110100daff01202010c0014a003274420b81),
    .INIT_4F(256'h0033021d001201ec0032cc0b03201100001a00209d00101c000380209c320b5c),
    .INIT_50(256'h014a00227c120b5c00d3ff0502020b81014a00208fa0101c00d2ff3270701100),
    .INIT_51(256'h0003800b01620b5c00021020f6020a60014b082f21e20b5c00daff0120420a63),
    .INIT_52(256'h00d2ff1d0ff20beb0033042f1152d0110032f02f01401002001a000b11720a66),
    .INIT_53(256'h00daff0b11920b3e014a000b01820beb00d3ff3483f2d011014a001f1ff01002),
    .INIT_54(256'h0009501f1ff202020250001d0ff20a5602fb272f115201bb014b082f014201b1),
    .INIT_55(256'h01490e2f014011000011000b11b201f700100c0b01a011000008403483f01010),
    .INIT_56(256'h036d573483f202020190011f1ff20b4c0131001d0ff20b810148082f11501010),
    .INIT_57(256'h0018ff2f115011000019ff2f014201f7036d610b11d0110001d1000b01c01014),
    .INIT_58(256'h0011020b0321d002036d673483f0b00200d5081f1ff20b810250001d0ff01014),
    .INIT_59(256'h01d1031d000010180250000b013202020018ff3677620b520019ff1d00032178),
    .INIT_5A(256'h0018ff1d0020101800004032771011000001501d001201f703ed743276f01100),
    .INIT_5B(256'h03ed6c20bb032178014008327751d00301410e1d0030b0020118013277320b81),
    .INIT_5C(256'h02500020bc501100001104227760101c00190b20bba202020118082277620b5c),
    .INIT_5D(256'h01b905209c320b81019818209d80101c00084020bd00110000095022776201f7),
    .INIT_5E(256'h0018ff1d0010300f0019ff0b03209001001102209d02b04e03ed7d20a00201b1),
    .INIT_5F(256'h014106227c10d00200381f030df09002000180208fa3219f025000327071d001),
    .INIT_60(256'h014106208dd2b40f014900208bf2b20f0141063678d20b120149001d00832190),
    .INIT_61(256'h036d8a0b0322b10f01d90b209a82b08f0011022089b2b04f014900208bf2b80f),
    .INIT_62(256'h025000050202d010001104208fa0101c03ad8c327072d01001d8141d001010e0),
    .INIT_63(256'h037001208bb220080250003679a2093a03ad8a1d0102090c01d808227c101002),
    .INIT_64(256'h00b40e209a81d00200b30d2089b0b00200b20c208e920216020e69208e32020d),
    .INIT_65(256'h01450e208fa1d003003403327070b0020005401d0012021f00ba0f0b0323219a),
    .INIT_66(256'h0007a0367a7010000036071d02020b120006a0227c12022801450e050203219a),
    .INIT_67(256'h01470e2089b20b1201470e208e92200801470e208e32093a01470e208bb2090c),
    .INIT_68(256'h000820327072b04f001e001d0012b80f001d000b0322b40f003703209a82b20f),
    .INIT_69(256'h032df31d0402d01001d603227c1010e0032dcb030df2b10f01d602208fa2b08f),
    .INIT_6A(256'h001a00208e92f032001900208e301001032e29208bb2d01001d604367b40101c),
    .INIT_6B(256'h032db71d0012089d01ce400b032208a1036db0209a8208c101cd302089b20928),
    .INIT_6C(256'h013a00227c12089b013900030df208cf0108f0208fa208d7009f0832707226cf),
    .INIT_6D(256'h001d00208d7208bb022dac208dd208bf013e0036017208cb011d011d08025000),
    .INIT_6E(256'h032dc10b032208cb01cd50209a82500000bf312089b2089d00be30208d3208d9),
    .INIT_6F(256'h011d01030df2089d013a00208fa208e10129f032707208cb0108e01d001208d5),
    .INIT_70(256'h003a032090c208bd02f91101008208c102f81020900208dd022dba227c125000),
    .INIT_71(256'h004a00367e5208c50140061d004250000140060b01e2089d00b01322008208cf),
    .INIT_72(256'h00bd30227ce0300f0250000504009001037000208fa2089d02fa12327c9208df),
    .INIT_73(256'h001a000b00e208bb001900209002500000b237030bf2089b00be31208fa20874),
    .INIT_74(256'h0108d0367e103008032dd8190010900201cf200b01f2089d001f002f03b208c5),
    .INIT_75(256'h022dd11d00220874011f010b0021400e013a00202451400e0129e02023c1400e),
    .INIT_76(256'h032de11d0030110001cf500b002010c000b23c2024e25000001f00327de2089b),
    .INIT_77(256'h011f010100201d01013a0020b1201e000139002025701f00010820327de20b6a),
    .INIT_78(256'h032de920922010a001cf300108225000001f002f01f20b98022dda2280f01c00),
    .INIT_79(256'h011f011d00801e000138003280001f000139001d00220b6a0118022200801100),
    .INIT_7A(256'h003a031d0202500002f9113280020b9802f8101d01001c00022de23280001d00),
    .INIT_7B(256'h004a002090003d7c0140060504003e3c014006208fa03f8100b013367f220b88),
    .INIT_7C(256'h00bd30367f905d030250001d04005e400370002280f05f0002fa120100203c3f),
    .INIT_7D(256'h0019000100220b88001800209002500000b237030bf20b9800be31208fa05c00),
    .INIT_7E(256'h032e01208fa03cff01cf203601703dfd001f001d08003e7f001a002280f03fff),
    .INIT_7F(256'h011f012280f05c00013a000100205d000129e02090005e800108d0030bf05f00),
    .INITP_00(256'hc3f2cee1726079514b01671fcdb6d419fda67100e10e44ab2d1739f8ece6b864),
    .INITP_01(256'h5d0bb3c8a6e126debb5f0f7b6bcae8760793972b63cd4fefedaf49b9e5994c29),
    .INITP_02(256'h1d898d889f1a08ab112e119f85cf51e3eb5c26a44d862897c69f13a3c82019a5),
    .INITP_03(256'h062b1aa609330a2fea32823a383e0c3210b02da8b5917b6ecd3cb78cea1d3988),
    .INITP_04(256'h613b92340c0983ba34afa1841a25d25e4713a50ec9363f2a11a5372b9c208bb1),
    .INITP_05(256'hbc9a221e0d3e5ffdcf04360b69819fae80071e1f160b848daa99ae051213a523),
    .INITP_06(256'hc50b27b0d92e05823402981610a931b638058ca20d172297e320162e04b5a53d),
    .INITP_07(256'h973cbbba9a0fab82133c2609059babbffda495ad3818a0b90d373235ab9551cc),
    .INITP_08(256'h18f689a0192a8c9a87b006b0b6ada747d1301e99a69e380e12b52dcfcd929a2b),
    .INITP_09(256'h3b1f9714a4192f3a2e8c3da2842c2f2ea5dd0cb1a9840d8e962431948a35fc6c),
    .INITP_0A(256'h9d92f917761c888a81161a1d91c3e531bf2fa8119cac8e368314033239b41497),
    .INITP_0B(256'h9d8212518a9504d334328094d026af8b49189937119dba5a3ce1983103fc88d7),
    .INITP_0C(256'ha4959a3822b1283632a0b9803aa1006a5dd3e7275b29603549a6193333aca007),
    .INITP_0D(256'h0cbc9a2a6516369f8dca86a38721872e7d8ef1a33930e8364e39433011003b2d),
    .INITP_0E(256'h99b0103dff1da73fca9f13b7914a3e0e0e0e862c33ec4b428581a38ab96c6f54),
    .INITP_0F(256'h1d930a82c4958484043983bcb8747de38d3f1ea61b5a5146b7042708e5388e55),
